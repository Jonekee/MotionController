Library IEEE;
use IEEE.std_logic_1164.all;

Entity SineLUTA is
	port(
	EANG : in std_logic_vector(3 downto 0);
	SINA : out std_logic_vector(17 downto 0);
	SINB : out std_logic_vector(17 downto 0)
	);
end SineLUTA;

Architecture DataFlow of SineLUTA is
begin
	With EANG Select SINA <=
	"000000000000000000" when "1011", --sin(0.00)
	"000110000111110111" when "1010", --sin(22.50)
	"001011010100000100" when "1110", --sin(45.00)
	"001110110010000010" when "1111", --sin(67.50)
	"001111111111111111" when "1101", --sin(90.00)
	"001110110010000010" when "1100", --sin(112.50)
	"001011010100000100" when "0100", --sin(135.00)
	"000110000111110111" when "0101", --sin(157.50)
	"000000000000000000" when "0111", --sin(180.00)
	"111001111000001001" when "0110", --sin(202.50)
	"110100101011111100" when "0010", --sin(225.00)
	"110001001101111110" when "0011", --sin(247.50)
	"110000000000000001" when "0001", --sin(270.00)
	"110001001101111110" when "0000", --sin(292.50)
	"110100101011111100" when "1000", --sin(315.00)
	"111001111000001001" when others; --sin(337.50)
	With EANG Select SINB <=
	"110010001001001110" when "1011", --sin(-120.00)
	"110000001000110010" when "1010", --sin(-97.50)
	"110000100010111011" when "1110", --sin(-75.00)
	"110011010011101000" when "1111", --sin(-52.50)
	"111000000000000001" when "1101", --sin(-30.00)
	"111101111010010110" when "1100", --sin(-7.50)
	"000100001001000001" when "0100", --sin(15.00)
	"001001101111010111" when "0101", --sin(37.50)
	"001101110110110010" when "0111", --sin(60.00)
	"001111110111001110" when "0110", --sin(82.50)
	"001111011101000101" when "0010", --sin(105.00)
	"001100101100011000" when "0011", --sin(127.50)
	"000111111111111111" when "0001", --sin(150.00)
	"000010000101101010" when "0000", --sin(172.50)
	"111011110110111111" when "1000", --sin(195.00)
	"110110010000101001" when others; --sin(217.50)
end DataFlow;